// Ejemplo: Hola mundo: holaMundoVerilog.v

module hello;
    initial
        $display ("Hola, mundo !!!");
endmodule