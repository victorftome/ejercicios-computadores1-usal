module ejer11;
	initial
	begin
		$display ("Decimal del numero %h : %d", 'h1FEA, 'h1FEA);
		$display ("Decimal del numero %b : %d", 7'b1000101, 7'b1000101);
		$display ("Octal del numero %d : %o", 1234, 1234);
		$display ("Hexadecimal del numero binario %b :%h", 7'b1010011, 7'b1010011);
	end
endmodule
